module led_module(
    input led_state,
    output led_out
);

assign led_out = led_state;

endmodule
